module xor_gate(a,b,xor_out);
    input a,b;
    output xor_out;
    assign xor_out= a^b;
endmodule
