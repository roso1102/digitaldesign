module not_gate(a,not_out);
    input a;
    output not_out;
    assign not_out= ~a;
endmodule