module buffer(a,buffer_out);
    input a;
    output buffer_out;
    assign buffer_out= a;
endmodule