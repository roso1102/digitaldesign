module or_gate(a,b,or_out);
    input a,b;
    output or_out;
    assign or_out= a | b;
endmodule